/*
Copyright by Henry Ko and Nicola Nicolici
Developed for the Digital Systems Design course (COE3DQ4)
Department of Electrical and Computer Engineering
McMaster University
Ontario, Canada
*/

`timescale 1ns/100ps
`default_nettype none

`include "define_state.h"

// This is the top module
// It connects the SRAM and VGA together
// It will first write RGB data of an image with 8x8 rectangles of size 40x30 pixels into the SRAM
// The VGA will then read the SRAM and display the image
module project (
		/////// board clocks                      ////////////
		input logic CLOCK_50_I,                   // 50 MHz clock

		/////// pushbuttons/switches              ////////////
		input logic[3:0] PUSH_BUTTON_I,           // pushbuttons
		input logic[17:0] SWITCH_I,               // toggle switches

		/////// VGA interface                     ////////////
		output logic VGA_CLOCK_O,                 // VGA clock
		output logic VGA_HSYNC_O,                 // VGA H_SYNC
		output logic VGA_VSYNC_O,                 // VGA V_SYNC
		output logic VGA_BLANK_O,                 // VGA BLANK
		output logic VGA_SYNC_O,                  // VGA SYNC
		output logic[9:0] VGA_RED_O,              // VGA red
		output logic[9:0] VGA_GREEN_O,            // VGA green
		output logic[9:0] VGA_BLUE_O,             // VGA blue
		
		/////// SRAM Interface                    ////////////
		inout wire[15:0] SRAM_DATA_IO,            // SRAM data bus 16 bits
		output logic[17:0] SRAM_ADDRESS_O,        // SRAM address bus 18 bits
		output logic SRAM_UB_N_O,                 // SRAM high-byte data mask 
		output logic SRAM_LB_N_O,                 // SRAM low-byte data mask 
		output logic SRAM_WE_N_O,                 // SRAM write enable
		output logic SRAM_CE_N_O,                 // SRAM chip enable
		output logic SRAM_OE_N_O                  // SRAM output logic enable
);

parameter NUM_ROW_RECTANGLE = 8,
		  NUM_COL_RECTANGLE = 8,
		  RECT_WIDTH = 40,
		  RECT_HEIGHT = 30,
		  VIEW_AREA_LEFT = 160,
		  VIEW_AREA_RIGHT = 480,
		  VIEW_AREA_TOP = 120,
		  VIEW_AREA_BOTTOM = 360;

parameter Y_OFFSET = 0, U_OFFSET = 18'd38400, V_OFFSET = 18'd57600, RGB_OFFSET = 18'd146944;

// Define the offset for Green and Blue data in the memory		
parameter RED_OFFSET = 18'd146944,
	  GREEN_EVEN_OFFSET = 18'd185344,
	  GREEN_ODD_OFFSET = 18'd204544,
	  BLUE_EVEN_OFFSET = 18'd223744,
	  BLUE_ODD_OFFSET = 18'd242944;

parameter U_21_CONSTANT = 32'd21, U_52_CONSTANT = 32'd52, U_159_CONSTANT = 32'd159;
parameter R_76284_CONSTANT = 32'd76284, R_25624_CONSTANT = 32'd25624, R_132251_CONSTANT = 32'd132251, R_104595_CONSTANT = 32'd104595, R_53281_CONSTANT = 32'd53281;

// Data counter for getting RGB data of a pixel
logic [17:0] data_counter;
state_top state;
logic done;

//keep track of whether or not we are working on an even collumn.
logic even_counter;

assign even_counter = ~data_counter[0];

logic [2:0] S_IDLE_WAIT;
// For Push button
logic [3:0] PB_pushed;

// For VGA
logic [9:0] VGA_red, VGA_green, VGA_blue;
logic [9:0] pixel_X_pos;
logic [9:0] pixel_Y_pos;

logic resetn;

// For SRAM
logic [17:0] SRAM_address;
logic [15:0] SRAM_write_data;
logic SRAM_we_n;
logic [15:0] SRAM_read_data;
logic [7:0] SRAM_read_high_byte, SRAM_read_low_byte;
logic SRAM_ready;

assign SRAM_read_high_byte = SRAM_read_data[15:8];
assign SRAM_read_low_byte = SRAM_read_data[7:0];

// For Colorspace conversion
logic [7:0] RED, GREEN, BLUE, Y_ODD, Y_EVEN, U_ODD, U_EVEN, V_ODD, V_EVEN, Y_multi_EVEN, U_multi_EVEN, V_multi_EVEN, Y_multi_ODD, U_multi_ODD, V_multi_ODD;

//logic [32:0]  

logic [31:0] U_21, U_52, U_159, V_21, V_52, V_159;

logic [63:0] R_result_EVEN, G_result_EVEN, B_result_EVEN, R_result_ODD, G_result_ODD, B_result_ODD;

logic [7:0] R_writable, G_writable, B_writable;

logic [8:0] U_N [7:0];
logic [8:0] V_N [7:0];

assign U_21 = U_N[5] + U_N[0];
assign U_52 = U_N[4] + U_N[1];
assign U_159 = U_N[3] + U_N[2];

assign V_21 = V_N[5] + V_N[0];
assign V_52 = V_N[4] + V_N[1];
assign V_159 = V_N[3] + V_N[2];

assign Y_multi_EVEN = Y_EVEN - 16;
assign U_multi_EVEN = U_EVEN - 128;
assign V_multi_EVEN = V_EVEN - 128;

assign Y_multi_ODD = Y_ODD - 16;
assign U_multi_ODD = U_ODD - 128;
assign V_multi_ODD = V_ODD - 128;

logic [31:0] mul0_op1, mul0_op2, mul0_result;
logic [31:0] mul1_op1, mul1_op2, mul1_result;
logic [31:0] mul2_op1, mul2_op2, mul2_result;

logic [2:0] rect_row_count;	// Number of rectangles in a row
logic [2:0] rect_col_count;	// Number of rectangles in a column
logic [5:0] rect_width_count;	// Width of each rectangle
logic [4:0] rect_height_count;	// Height of each rectangle
logic [2:0] color;

logic [15:0] VGA_sram_data [2:0];

logic [7:0] Red_buf, G2_buf, B2_buf;

logic RED_second_word;

assign resetn = ~SWITCH_I[17] && SRAM_ready;

// Push Button unit
PB_Controller PB_unit (
	.Clock_50(CLOCK_50_I),
	.Resetn(resetn),
	.PB_signal(PUSH_BUTTON_I),	
	.PB_pushed(PB_pushed)
);

// SRAM unit
SRAM_Controller SRAM_unit (
	.Clock_50(CLOCK_50_I),
	.Resetn(~SWITCH_I[17]),
	.SRAM_address(SRAM_address),
	.SRAM_write_data(SRAM_write_data),
	.SRAM_we_n(SRAM_we_n),
	.SRAM_read_data(SRAM_read_data),		
	.SRAM_ready(SRAM_ready),
		
	// To the SRAM pins
	.SRAM_DATA_IO(SRAM_DATA_IO),
	.SRAM_ADDRESS_O(SRAM_ADDRESS_O),
	.SRAM_UB_N_O(SRAM_UB_N_O),
	.SRAM_LB_N_O(SRAM_LB_N_O),
	.SRAM_WE_N_O(SRAM_WE_N_O),
	.SRAM_CE_N_O(SRAM_CE_N_O),
	.SRAM_OE_N_O(SRAM_OE_N_O)
);

// VGA unit
VGA_Controller VGA_unit(
	.Clock(CLOCK_50_I),
	.Resetn(resetn),

	.iRed(VGA_red),
	.iGreen(VGA_green),
	.iBlue(VGA_blue),
	.oCoord_X(pixel_X_pos),
	.oCoord_Y(pixel_Y_pos),
	
	//	VGA Side
	.oVGA_R(VGA_RED_O),
	.oVGA_G(VGA_GREEN_O),
	.oVGA_B(VGA_BLUE_O),
	.oVGA_H_SYNC(VGA_HSYNC_O),
	.oVGA_V_SYNC(VGA_VSYNC_O),
	.oVGA_SYNC(VGA_SYNC_O),
	.oVGA_BLANK(VGA_BLANK_O),
	.oVGA_CLOCK(VGA_CLOCK_O)
);

milestone1_multiplier mul0 (
	.Resetn(resetn),
	.value00(mul0_op1),
	.value01(mul0_op2),
	.select(1'b0),
	.result(mul0_result)
);

milestone1_multiplier mul1 (
	.Resetn(resetn),
	.value00(mul1_op1),
	.value01(mul1_op2),
	.select(1'b0),
	.result(mul1_result)
);

milestone1_multiplier mul2 (
	.Resetn(resetn),
	.value00(mul2_op1),
	.value01(mul2_op2),
	.select(1'b0),
	.result(mul2_result)
);


// Each rectangle will have different color
assign color = rect_col_count + rect_row_count;

always_ff @ (posedge CLOCK_50_I or negedge resetn) begin
	if (resetn == 1'b0) begin
		state <= S_IDLE_TOP;
		S_IDLE_WAIT <= 2'b00;
		rect_row_count <= 3'd0;
		rect_col_count <= 3'd0;
		rect_width_count <= 6'd0;
		rect_height_count <= 5'd0;
		
		VGA_red <= 10'd0;
		VGA_green <= 10'd0;
		VGA_blue <= 10'd0;				
		
		SRAM_we_n <= 1'b1;
		SRAM_write_data <= 16'd0;
		SRAM_address <= 18'd0;
		
		data_counter <= 18'd0;
		RED_second_word <= 1'b0;

		Y_ODD <= 1'b0;
		Y_EVEN <= 1'b0;
		U_ODD <= 1'b0;
		U_EVEN <= 1'b0;
		V_ODD <= 1'b0;
		V_EVEN <= 1'b0;

		U_N[0] <= 1'b0;
		U_N[1] <= 1'b0;
		U_N[2] <= 1'b0;
		U_N[3] <= 1'b0;
		U_N[4] <= 1'b0;
		U_N[5] <= 1'b0;
		U_N[6] <= 1'b0;
		U_N[7] <= 1'b0;

		V_N[0] <= 1'b0;
		V_N[1] <= 1'b0;
		V_N[2] <= 1'b0;
		V_N[3] <= 1'b0;
		V_N[4] <= 1'b0;
		V_N[5] <= 1'b0;
		V_N[6] <= 1'b0;
		V_N[7] <= 1'b0;

	end else begin
		case (state)
		S_IDLE_TOP: begin
			S_IDLE_WAIT <= S_IDLE_WAIT + 1'b1;
			if (S_IDLE_WAIT == 2'b1) begin
				S_IDLE_WAIT <= 1'b0;
				state <= S_READ_U_0;
				SRAM_address <= data_counter + U_OFFSET;
			end
			done <= 1'b1;
		end

		S_READ_U_0: begin
			state <= S_READ_U_1;
			SRAM_address <= data_counter + U_OFFSET + 1; 
		end

		S_READ_U_1: begin
			state <= S_READ_V_0;
			SRAM_address <= data_counter + V_OFFSET; 
		end

		S_READ_V_0: begin
			SRAM_address <= data_counter + V_OFFSET + 1; 
			U_EVEN <= SRAM_read_high_byte;
			U_N[0] <= SRAM_read_high_byte;
			U_N[1] <= SRAM_read_high_byte;
			U_N[2] <= SRAM_read_high_byte;
			U_N[3] <= SRAM_read_low_byte;
			state <= S_READ_V_1;

		end
		
		S_READ_V_1: begin
			SRAM_address <= data_counter + Y_OFFSET;
			U_N[4] <= SRAM_read_high_byte;
			U_N[5] <= SRAM_read_low_byte;
			state <= S_READ_Y;
		end

		S_READ_Y: begin
			V_EVEN <= SRAM_read_high_byte;
			V_N[0] <= SRAM_read_high_byte;
			V_N[1] <= SRAM_read_high_byte;
			V_N[2] <= SRAM_read_high_byte;
			V_N[3] <= SRAM_read_low_byte;
			state <= S_START_ROW;
		end
		S_START_ROW: begin
			V_N[4] <= SRAM_read_high_byte;
			V_N[5] <= SRAM_read_low_byte;
			
			state <= S_CALC_U;
		end
		S_CALC_U: begin


			mul0_op1 <= U_21;
			mul0_op2 <= U_21_CONSTANT;
			mul1_op1 <= U_52;
			mul1_op2 <= U_52_CONSTANT;
			mul2_op1 <= U_159;
			mul2_op2 <= U_159_CONSTANT;

			state <= S_CALC_V;
		end

		S_CALC_V: begin

			U_ODD <= mul0_result - mul1_result + mul2_result + 128;

			mul0_op1 <= V_21;
			mul0_op2 <= U_21_CONSTANT;
			mul1_op1 <= V_52;
			mul1_op2 <= U_52_CONSTANT;
			mul2_op1 <= V_159;
			mul2_op2 <= U_159_CONSTANT;

			//load Y
			Y_EVEN <= SRAM_read_high_byte;
			Y_ODD <= SRAM_read_low_byte;
			
			state <= S_CALC_R00;
		end

		S_CALC_R00: begin
			V_ODD <= mul0_result - mul1_result + mul2_result + 128;

			mul0_op1 <= Y_multi_EVEN;
			mul0_op2 <= R_76284_CONSTANT;

			mul1_op1 <= U_multi_EVEN;
			mul1_op2 <= R_25624_CONSTANT;

			mul2_op1 <= V_multi_EVEN;
			mul2_op2 <= R_104595_CONSTANT;

			state <= S_CALC_R01;
		end

		S_CALC_R01: begin

			R_result_EVEN <= mul0_result + mul2_result;
			G_result_EVEN <= mul0_result - mul1_result;
			B_result_EVEN <= mul0_result;

			mul0_op1 <= 0;
			mul0_op2 <= 0;

			mul1_op2 <= R_132251_CONSTANT;

			mul2_op2 <= R_53281_CONSTANT;
			
			state <= S_CALC_R10;
		end


		S_CALC_R10: begin

			G_result_EVEN <= G_result_EVEN - mul2_result;
			B_result_EVEN <= B_result_EVEN + mul1_result;

			mul0_op1 <= Y_multi_ODD;
			mul0_op2 <= R_76284_CONSTANT;

			mul1_op1 <= U_multi_ODD;
			mul1_op2 <= R_25624_CONSTANT;

			mul2_op1 <= V_multi_ODD;
			mul2_op2 <= R_104595_CONSTANT;
			
			state <= S_CALC_R11;
		end

		S_CALC_R11: begin

			R_result_ODD <= mul0_result + mul2_result;
			G_result_ODD <= mul0_result - mul1_result;
			B_result_ODD <= mul0_result;

			mul0_op1 <= 0;
			mul0_op2 <= 0;

			mul1_op2 <= R_132251_CONSTANT;

			mul2_op2 <= R_53281_CONSTANT;
			
			state <= S_IDLE_TOP;
		end

		default: state <= S_IDLE_TOP;
		endcase
	end
end

endmodule
